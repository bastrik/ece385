// The datapath module should handle 

module datapath(
);

endmodule