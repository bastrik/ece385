// Arithmetic logic unit

module ALU (input logic [15:0] A, B,
            input logic [1:0] select,
            output logic [15:0] out);

always_comb
begin

	case (select)
	       // ADD
	       2'b00:
		       out = A + B;
	       // AND
	       2'b01:
		       out = A & B;
	       // NOT A
	       2'b10:
		       out = ~A;
	       // PASS A
	       2'b11:
		       out = A;
       endcase
end

endmodule
